0 1 0
1 1 1
2 1 2
3 1 3
4 1 4
5 1 5
6 1 6
7 1 7
8 1 8
9 1 9
10 1 10
11 1 11
12 1 12
13 1 13
14 1 14
15 1 15
16 1 16
17 1 17
18 1 18
19 1 19
20 1 20
21 1 21
22 1 22
23 1 23
24 1 24
25 1 25
26 1 26
27 1 27
28 1 28
29 1 29
30 1 30
31 1 31
32 1 32
33 1 33
34 1 34
35 1 35
36 3 36
37 3 37
38 3 38
39 3 39
40 3 40
41 3 41
42 3 42
43 0 5 44 43
44 0 5 45 43
45 0 5 46 43
46 0 5 47 43
47 0 5 48 43
48 0 5 49 43
49 0 5 50 43
50 0 5 51 43
51 0 5 52 43
52 0 5 53 43
53 0 5 54 43
54 0 5 55 43
55 0 5 56 43
56 0 5 57 43
57 0 5 58 43
58 0 5 59 43
59 0 5 60 43
60 0 5 61 43
61 0 6 62 44 1
62 0 3 63 2 45
63 0 3 64 4 45
64 0 6 65 46 5
65 0 6 66 48 9
66 0 6 67 50 13
67 0 6 68 52 17
68 0 6 69 54 21
69 0 6 70 56 25
70 0 6 71 58 29
71 0 6 72 60 33
72 0 3 73 6 47
73 0 3 74 8 47
74 0 3 75 10 49
75 0 3 76 12 49
76 0 3 77 14 51
77 0 3 78 16 51
78 0 3 79 18 53
79 0 3 80 20 53
80 0 3 81 22 55
81 0 3 82 24 55
82 0 3 83 26 57
83 0 3 84 28 57
84 0 3 85 30 59
85 0 3 86 32 59
86 0 3 87 34 61
87 0 3 88 35 61
88 0 1 62 65
89 0 5 90 43
90 0 5 91 43
91 0 5 92 43
92 0 5 93 43
93 0 6 94 90 93
94 0 6 95 62 92
95 0 6 96 94 95
96 0 5 97 43
97 0 5 98 43
98 0 6 99 90 98
99 0 6 100 65 97
100 0 6 101 99 100
101 0 5 102 43
102 0 5 103 43
103 0 6 104 90 103
104 0 6 105 66 102
105 0 6 106 104 105
106 0 5 107 43
107 0 5 108 43
108 0 6 109 90 108
109 0 6 110 67 107
110 0 6 111 109 110
111 0 5 112 43
112 0 5 113 43
113 0 6 114 90 113
114 0 6 115 68 112
115 0 6 116 114 115
116 0 5 117 43
117 0 5 118 43
118 0 6 119 90 118
119 0 6 120 69 117
120 0 6 121 119 120
121 0 6 122 0 91
122 0 5 123 43
123 0 5 124 43
124 0 6 125 90 124
125 0 6 126 70 123
126 0 6 127 125 126
127 0 6 128 91 3
128 0 5 129 43
129 0 5 130 43
130 0 6 131 90 130
131 0 6 132 71 129
132 0 6 133 131 132
133 0 6 134 91 7
134 0 5 135 43
135 0 5 136 43
136 0 6 137 90 136
137 0 6 138 72 135
138 0 6 139 137 138
139 0 6 140 91 11
140 0 6 141 91 15
141 0 6 142 91 19
142 0 6 143 91 23
143 0 6 144 91 27
144 0 6 145 91 31
145 0 6 146 96 63
146 0 6 147 96 64
147 0 6 148 101 73
148 0 6 149 106 75
149 0 6 150 111 77
150 0 6 151 116 79
151 0 6 152 121 81
152 0 6 153 127 83
153 0 6 154 133 85
154 0 6 155 139 87
155 0 6 156 101 74
156 0 6 157 106 76
157 0 6 158 111 78
158 0 6 159 116 80
159 0 6 160 121 82
160 0 6 161 127 84
161 0 6 162 133 86
162 0 6 163 139 88
163 0 1 146 148
164 0 5 165 43
165 0 5 166 43
166 0 5 167 43
167 0 5 168 43
168 0 5 169 43
169 0 5 170 43
170 0 5 171 43
171 0 5 172 43
172 0 5 173 43
173 0 5 174 43
174 0 5 175 43
175 0 5 176 43
176 0 5 177 43
177 0 6 178 174 177
178 0 6 179 146 176
179 0 6 180 178 179
180 0 5 181 43
181 0 5 182 43
182 0 6 183 174 182
183 0 6 184 148 181
184 0 6 185 183 184
185 0 5 186 43
186 0 5 187 43
187 0 6 188 174 187
188 0 6 189 149 186
189 0 6 190 188 189
190 0 5 191 43
191 0 5 192 43
192 0 6 193 174 192
193 0 6 194 150 191
194 0 6 195 193 194
195 0 6 196 2 175
196 0 5 197 43
197 0 5 198 43
198 0 6 199 174 198
199 0 6 200 151 197
200 0 6 201 199 200
201 0 6 202 175 6
202 0 5 203 43
203 0 5 204 43
204 0 6 205 174 204
205 0 6 206 152 203
206 0 6 207 205 206
207 0 6 208 175 10
208 0 5 209 43
209 0 5 210 43
210 0 6 211 174 210
211 0 6 212 153 209
212 0 6 213 211 212
213 0 6 214 175 14
214 0 5 215 43
215 0 5 216 43
216 0 6 217 174 216
217 0 6 218 154 215
218 0 6 219 217 218
219 0 6 220 175 18
220 0 5 221 43
221 0 5 222 43
222 0 6 223 174 222
223 0 6 224 155 221
224 0 6 225 223 224
225 0 6 226 175 22
226 0 6 227 175 26
227 0 6 228 175 30
228 0 6 229 175 34
229 0 6 230 180 165
230 0 6 231 185 166
231 0 6 232 190 167
232 0 6 233 195 168
233 0 6 234 201 169
234 0 6 235 207 170
235 0 6 236 213 171
236 0 6 237 219 172
237 0 6 238 225 173
238 0 1 230 231
239 0 5 240 43
240 0 6 241 4 240
241 0 6 242 240 8
242 0 6 243 240 12
243 0 6 244 240 16
244 0 6 245 240 20
245 0 6 246 240 24
246 0 6 247 240 28
247 0 6 248 240 32
248 0 6 249 240 35
249 0 6 250 1 122
250 0 6 251 128 202
251 0 6 252 134 208
252 0 6 253 140 214
253 0 6 254 141 220
254 0 6 255 142 226
255 0 6 256 143 227
256 0 6 257 144 228
257 0 6 258 145 229
258 0 5 259 43
259 0 1 251 252
260 0 5 261 43
261 0 5 262 43
262 0 5 263 43
263 0 5 264 43
264 0 6 265 252 261
265 0 6 266 252 253
266 0 6 267 254 253
267 0 6 268 252 253
268 0 5 36 43
269 0 5 37 43
270 0 5 38 43
271 0 3 39 259 260
272 0 6 40 251 252
273 0 6 41 251 252
274 0 6 42 251 265

0 1 0
1 1 1
2 1 2
3 1 3
4 1 4
5 3 5
6 3 6
7 0 6 7 0 2
8 0 6 8 2 3
9 0 6 9 1 8
10 0 6 10 8 4
11 0 6 5 7 9
12 0 6 6 9 10
